`timescale 1ns/1ps

module tb_layer_one_trained;

    // =========================================================
    // Actual trained weights from layer_0_weights.mem
    // Actual thresholds from layer_1_thresholds.mem
    // Real MNIST test images from mnist_binary_verifying.ubin
    // =========================================================

    // Trained weights (same for all tests)
    reg [71:0] TRAINED_WEIGHTS = 72'b000001100000011100000011100001101000110110001111111110000111100011101010;

    // Image 0: MNIST label=5, active outputs=883/1568
    reg [783:0]  PIXELS_0   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001111111100000000000000000001111111111000000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000011111111111100000000000000000111111111111000000000000000000001100011110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000011111000000000000000000001111111100000000000000000111111111100000000000000111111111111100000000000000111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_0 = 1568'b00000000000000000000110000000001111100000000110000000000000000000000000000110000000000000111111000000000000011000000000000000000000011110000000111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111011111111111101111111111111011111111111111011111111111111111101111111111111101111111111111011111111110001111111000111111111111111111111111111111111111111111111111111111111111111111111101111111111000111111111110111111111111101111111111111100111111111111110010011111111111110111111111111001111111111000011111100011011111111111111111111111111111111111111111111111111111111111111111110111111111100111111111111011111111111110111111111111110011111111111111111011111111111111111111111111101111111111100011111111011111111111111111111111111111111111110000000000000000001111000000000111110000000011000000000000010000000000000011111100000000011111100000000000001000000000001100000000011111000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000111111000000001100000000000011000000000000111111100000000011111110000000000001100000000000111000000011111110000111111111000000000000000000000000000000000000000000000000000000000000000111100000000111111000000001100000000000001100000000000011111110000000001111110000000000001100000000000011000000000111110000001111111000000000000000000000000000000001111111111111111111101111111111111110111111111111111111111110111111111111110111111111111111111011111111111110111111111111101111111111011111111100111111111111111111111111111111111111111111111111111;

    // Image 1: MNIST label=3, active outputs=869/1568
    reg [783:0]  PIXELS_1   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000111111111111000000000000000111110001111100000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000111111100000000000000000000111111110000000000000000000111111110000000000000000000110000000000000000000000001111000000000000000000000001100000000000000000000000001100000000000000000000000000111000000000000000000000000001111111111100000000000000000011111111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_1 = 1568'b00000000000000000000000000000000011111110000001000000000000010000000000000001000000000000011110000000001100000000001100000000000100000000000000111111000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110110011111111111111111111110111111111111111111111111111100011111111110111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111110001000111111101111111111111011111111111111111111111111110000111111111011111111111011111111111101111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111001110111111111111111111111101111111111111111111111111111000111111111111111111111111111111111111111111111111111000011111111111111111111111111111111110000000000000000000011111000000001111110000000110000000000001100000000000001100000000000001111000000001110000000000110000000000011000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000001111111000000111000000000001100000000000001110000000000011111000000001111110000000111000000000011100000000000011111100000000000111000000000000000000000000000000000000000000000000000001111100000001011111000000001000000000000110000000000000110000000000000111100000000111110000000001000000000001100000000000001111110000000000011000000000000000000001111111111111111111111111111111111111100111111111111111111111111111111111111011111111111111000111111111111101111111111111111111111111111111111110000011111111111110111111111111111111111111111111111;

    // Image 2: MNIST label=5, active outputs=876/1568
    reg [783:0]  PIXELS_2   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111110000000000000011111000000001100000000000011100000000000011000000000011100000000000000100000000011000000000000000010000000011000000000000000000000000001100000000000000110000000000110000000000000111000000000011100000000001111100000000000111000000111110110000000000001111111111100001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000011110000000000000000001111111110000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_2 = 1568'b00000000000000000000000000000000011111000000011110011000000100000001000100000000000000000000111000001100111100000001111000010000000000000000000001111100000000110000000000000000000000000000000000001111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111101111111000001111111111111111111111111111110111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111011111011111011111111011101111111111111011111110111111000000110111111111111101111111111111011111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111110111111111111111111111011111110000111111111111111111111111111111101111111100111111111111111111111111111111111110000000000000000000000000000000011111110000001110000100000110000000000011000000110000100000011100000111111100000000000000010000000000001100000001111110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000001111000110000111000000100001000000010000110000011100000111111101100000000000011000000000111110000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000111000010000001000000000001000000000000011000001100000011111111000000000000010000000000000110000000111111000000000000000000000000000000001111111111111111111111111111111111000011111110111111111111111111111111111111111111111101111111011111101101110111111111111111111111111111111111111101111111111111111111111111111111111111111111111111;

    // Image 3: MNIST label=0, active outputs=870/1568
    reg [783:0]  PIXELS_3   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111100000000000000001110000000111000000000000011100000000001100000000000011000000000000110000000000011000000000000110000000000011000000000000011000000000001100000000000011100000000001100000000000001100000000000110000000000011100000000000010000000000011100000000000001000000000001100000000000000000000000000100000000000000111000010101100000000000000011100111111100000000000000001110111111000000000000000000011111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_3 = 1568'b00000000000000000000000000000000000111110000000111000010000011000000000010000000100000100000010000000000001100000000001100000001111111100000000110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000011111111011111011111111111111111110111111111111111111111111111111111111111111111111111111011001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111101111101111110111111011111011111100111100111111011111111111101111111111110111111101100111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111110111111111111111111111111111111111111110000000000000000000000000000000000111111000000111000000000011000001100001100000010000011000001100000000000110000001000111000000111111100000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000111100011000001100000110000110000011000011000001110000110000111000001101111100000011111110000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000001100011000000100000000000000000000100001000000010000000000011000001100000100000001011110000000001110000000000000000000000000000000000001111111111111111111111111111111111100000111111111111101111111111111111111111111111111111111111101111101111111111111111111111111110001111111111101111111111111111111111111111111111111111111111111111;

    // Image 4: MNIST label=0, active outputs=851/1568
    reg [783:0]  PIXELS_4   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011111100000000000000000000011111110000000000000000000011111111100000000000000000001111101111000000000000000001111000001100000000000000001111000000110000000000000000111000000011000000000000000111100000001100000000000000011100000000110000000000000011100000000011000000000000001110000000001100000000000000110000000000110000000000000011000000000011000000000000000100000000001100000000000000011100000001110000000000000000111000000110000000000000000011111111111000000000000000000111111100100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_4 = 1568'b00000000000000000000000000000000001111000000001111110000000011000010000001100000000000011000000000001100000000000000000000000000011000100000000011111000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110011111111111100011111111110111011111111011110111111110111101111111011111011111111111111111111110111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111100000111111110011101111111100111011111110011110111111101111101111111011111011111111011110111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111110011111111111011111111111110111111111111011111111111110111111111111111111111111111101111111111111100011111111111111111111111111111111110000000000000000000001000000000001111000000000111011000000001100000000000110000100000001100001000000110000010000000100000100000001100011000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000111000000000011111100000001110011000000011000110000001110001100000011000011000000110000110000000110111100000001111110000000000111000000000000000000000000000000000000000000000000000000000000000000011100000000001111100000000101010000000000100100000001000001000000011000010000000010000000000000110001000000000111110000000000011000000000000000000001111111111111111111111111111111111010111111111111110111111111111111111111111111111111111101111111111110111111111111111111111111111011111111111111000101111111111111111111111111111111111111111111111;

    // Image 5: MNIST label=1, active outputs=823/1568
    reg [783:0]  PIXELS_5   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000001000000000000000000000000001100000000000000000000000001100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_5 = 1568'b00000000000000000000000000000000000111000000000001100000000000100000000000001000000000000110000000000001000000000000110000000000001000000000000001000000000001000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011111111111111111111111111011111111111101111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111101111111111110111111111111001111111111110111111111111001111111111110111111111111101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111111111011111111111101111111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000110000000000011100000000000110000000000011000000000000110000000000011000000000000110000000000011000000000000100000000000001000000000000110000000000000000000000000000000000000000000000000000000000000000000000000010000000000001100000000000111000000000001100000000000111000000000001100000000000111000000000011100000000000010000000000001100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000001010000000000010000000000000110000000000000000000000000000000000001111111111111111111111111111111111111011111111111110111111111111111111111111111111111111111011111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111;

    // Image 6: MNIST label=8, active outputs=863/1568
    reg [783:0]  PIXELS_6   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000011101100000000000000000000001100110000000000000000000001100011000000000000000000001100001000000000000000000000110000100000000000000000000011000110000000000000000000001100010000000000000000000000011111000000000000000000000000011110000000000000000000000001101000000000000000000000001100110000000000000000000000100001000000000000000000000110000100000000000000000000010000010000000000000000000011000011000000000000000000001100011000000000000000000000001011000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_6 = 1568'b00000000000000000000000000000000001110000000000110000000000010000000000000001100000000000111000000000000011000000000010110000000001100000000000010101000000000001000000000000000000000000000000000001111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111101001111111110011111111111101111111111111110011111111111100111111111110111111111111101101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001100000000001111000000000011100000000001100000000000010110000000000001100000000000110000000000001010000000000110110000000001011000000000001100000000000000000000000000000000000000000000000000000000000000000000001100000000000111000000000011110000000000101100000000011111000000000011100000000000011100000000001101000000000110110000000000111100000000000110000000000000000000000000000000000000000000000000000000100000000000011000000000000110000000000100000000000001100000000000001110000000000001100000000000001000000000001001000000000011100000000000010000000000000000000001111111111111111111111111111111111110111111111111101111111111111011111111110111111111111110111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111;

    // Image 7: MNIST label=4, active outputs=842/1568
    reg [783:0]  PIXELS_7   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000001111111100000000000000000000001111111110000000000000000000011111111100000000000000000001110011110000000000000000000110000110000000000000000000111000110000000000000000000011000011000000000000000000011000011000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_7 = 1568'b00000000000000000000000000000000000011000000000011100000000000110000000001111000000000000001110000000000000000000000100100000000010000000000001100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111101111111111111111111111111111111111111100111111111111111011111111110110111111111111011111111110111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111111111111111111111100001111111111100100111111111011011111111101101111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111101111111111111111111111111000111111111110110111111111101111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000110000000000011100000000001110000000000011000000000111101000000000000110000000001100000000000010010000000001100000000000110000000000001100000000000000000000000000000000000000000000000000000000000000000000000000010000000000001100000000000111000000011001100000000011111100000000011111000000000110110000000011111000000001110000000000111000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000001111100000000010111100000000010000000000000000100000000000000000000001100000000000000000000000000000000000001111111111111111111111111111111111111011111111111110111111111111111111111110111111111111111100111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

    // Image 8: MNIST label=3, active outputs=845/1568
    reg [783:0]  PIXELS_8   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111000000000000000000001111111100000000000000000001111111110000000000000000001111110000000000000000000000111100000000000000000000000011110000000000000000000000000111110000000000000000000000011111110000000000000000000000111111110000000000000000000001111111000000000000000000011111111100000000000000000001111111100000000000000000001111110000000000000000000001111100001000000000000000000111100000111000000000000000011111111111100000000000000000111111111110000000000000000001111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_8 = 1568'b00000000000000000000111100000000011100000000011100000000000000000000000000011110000000000001110000000011000000000001100110000000000111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100111111111100001111111110111111111111100111111111111110011111111111100011111111110011111111111011111111111110000011111111110001111111111111111111111111111111111111111111111111111111111111111111110011111111110000111111111001111111111110011111111111111001111111111100001111111111001111111111001111111111111000000111111111000111111111111111111111111111111111111111111111111111111111111111111111011111111111000111111111100111111111111101111111111111100111111111110000111111111101111111111110111111111111100000111111111110111111111111111111111111111111111110000000000000000000011100000000011110000000001110000000000001010000000000001111000000000010110000000001100000000000110011100000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000001111100000000111100000000001111000000000011111100000000011111000000001111100000000111001100000001111111000000001111110000000000000000000000000000000000000000000000000000000000000000001110000000000111100000000111100000000000111000000000001111100000000001111000000000111100000000011000100000000111111100000000111110000000000000000000000000000000001111111111111111111110011111111110110111111111111111111111111011111111111111001111111111110001111111111111111111111111110111111111100010111111111101101111111111111111111111111111111111111111111111;

    // Image 9: MNIST label=4, active outputs=860/1568
    reg [783:0]  PIXELS_9   = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001111111111110000000000000111111111111111100000000000001111000011111110000000000000110000000111110000000000000111000000111100000000000000011000000011100000000000000001000000011100000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_9 = 1568'b00000000000000000000000000000000001110000000000010000000000001000000000000010000000000011111111100000000000000000010000110000000000001000000000001100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110111000111111111110111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111110011111111111111111111111110011111111111001100011111100111001111111011100111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111001111111111101110001111110111101111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001100000000000111000000000001100000000000110000000000011011110000001111111100000010000100000001100011000000000001100000000000110000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000011000000000001110000000000011000000001101111110000001111111110000011000111000000110011100000000001100000000000111000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000111110000000111111110000010100001000000010001100000000000000000000000010000000000000000000000000000000000001111111111111111111111111111111111110111111111111101111111111111111111111111111111111111111100011111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111;

    // DUT signals
    reg clk, rst_n;
    reg [2:0] state;
    reg [783:0]  pixels;
    reg [71:0]   weights;
    wire [1567:0] layer_one_out;
    wire done;

    integer errors = 0, total_checks = 0;

    layer_one dut (
        .clk(clk), .rst_n(rst_n), .state(state),
        .pixels(pixels), .weights(weights),
        .layer_one_out(layer_one_out), .done(done)
    );

    localparam [2:0] s_LAYER_1 = 3'b010;

    initial begin clk = 0; forever #5 clk = ~clk; end

    function integer out_idx;
        input integer k, r, c;
        begin out_idx = k*196 + r*14 + c; end
    endfunction

    task run_test;
        input [783:0]  pix;
        input [1567:0] expected;
        input integer  img_idx;
        input integer  label;
        integer k, r, c, idx, mismatches;
        begin
            mismatches = 0;
            rst_n = 0; state = 3'b000;
            pixels = pix; weights = TRAINED_WEIGHTS;
            #20; rst_n = 1;
            #20; state = s_LAYER_1;
            wait(done == 1);
            #100;

            for (k = 0; k < 8; k = k + 1)
                for (r = 0; r < 14; r = r + 1)
                    for (c = 0; c < 14; c = c + 1) begin
                        idx = out_idx(k, r, c);
                        total_checks = total_checks + 1;
                        if (layer_one_out[idx] !== expected[idx]) begin
                            mismatches = mismatches + 1;
                            errors = errors + 1;
                        end
                    end

            if (mismatches == 0)
                $display("PASS  image=%0d  label=%0d", img_idx, label);
            else
                $display("FAIL  image=%0d  label=%0d  mismatches=%0d/1568", img_idx, label, mismatches);
        end
    endtask

    initial begin
        $dumpfile("layer_one_trained.vcd");
        $dumpvars(0, tb_layer_one_trained);

        $display("\n====================================================");
        $display("Layer One vs Trained Model - Real MNIST Test");
        $display("Weights: actual trained weights from layer_0_weights.mem");
        $display("Images:  real MNIST from mnist_binary_verifying.ubin");
        $display("Testing 10 images");
        $display("====================================================\n");

        run_test(PIXELS_0, EXPECTED_0, 0, 5);
        run_test(PIXELS_1, EXPECTED_1, 1, 3);
        run_test(PIXELS_2, EXPECTED_2, 2, 5);
        run_test(PIXELS_3, EXPECTED_3, 3, 0);
        run_test(PIXELS_4, EXPECTED_4, 4, 0);
        run_test(PIXELS_5, EXPECTED_5, 5, 1);
        run_test(PIXELS_6, EXPECTED_6, 6, 8);
        run_test(PIXELS_7, EXPECTED_7, 7, 4);
        run_test(PIXELS_8, EXPECTED_8, 8, 3);
        run_test(PIXELS_9, EXPECTED_9, 9, 4);

        $display("\n====================================================");
        if (errors == 0)
            $display("ALL 10 TESTS PASSED (%0d checks)", total_checks);
        else
            $display("FAILED: %0d errors / %0d checks", errors, total_checks);
        $display("====================================================\n");
        #50; $finish;
    end

    initial begin #200000000; $display("TIMEOUT"); $finish; end

endmodule
