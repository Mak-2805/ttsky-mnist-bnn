`timescale 1ns/1ps

// Define state_t here — avoids compiling fsm.sv which crashes icarus 10.2
// (fsm.sv uses always_ff/always_comb which trigger an assertion bug).
// layer_two.sv accepts the port connection because state_t is logic [2:0].
typedef enum logic [2:0] {
    s_IDLE    = 3'b000,
    s_LOAD    = 3'b001,
    s_LAYER_1 = 3'b010,
    s_LAYER_2 = 3'b011,
    s_LAYER_3 = 3'b100
} state_t;

module tb_layer_two;

    // ================================================================
    // Weights — packed as logic [2:0][2:0][7:0]
    //   bits [3:0] at each position = filter weights 3..0
    //   bits [7:4] unused (zero)
    //   Derived from layer_3_weights.mem via majority vote
    // ================================================================
    logic [2:0][2:0][7:0] TRAINED_WEIGHTS = 72'b000011000000101000001000000011010000110100001100000001110000111100001111;

    // ================================================================
    // Per-test pixel inputs and expected outputs
    //   pixels  : logic [13:0][13:0][7:0]  — 14x14 × 8-ch feature map
    //   expected: logic [3:0][6:0][6:0]    — 4 filters × 7x7
    // ================================================================
    // Image 0: label=5, active outputs=114/196
    logic [13:0][13:0][7:0] PIXELS_0   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011110011111100011111001011100010111000101110001011100010111000101110001011100010111000101110001111110011111111111111111110011111111111101110100011100010111000101110001011100010111000101110001011100011111101111001111000001110101011101110111011101110111010101110001011100010111000101110001011100010111000101110001011100110000111101110100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001000001111111111111111000011110010111100101111001011110010111000101110001011100010111000101110001011100010111000101110111000001111100111111111111111111111111111111111111111110000111000101110001011100010111000101110001011100010111000101110001011101110101011101010111011101110000011111011110111101010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011110110001011001110101011100010111000101110001011100010111000101110001011100010111100111111001111110001111100111001111000101110111010101110001011100010111000101110001011100011111100011111000111111011111111110001111000001110000011101010111011101010111000101110001011100010111000101110101000101110000011100010111011101110111011101010111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_0 = 196'b0111000111110011111000111111011111111111111111110111111111111111111111111111111111111111111111111100111000000000001110000000000000000000000000000001111111001110000111100001110001110000010000000000;

    // Image 1: label=3, active outputs=102/196
    logic [13:0][13:0][7:0] PIXELS_1   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101111001011110010111100101111001011100010111000101110001011100010111000101110001011100010111000111111001111111111111111111111111111111111111111011110100011100010111000101110001011100010111000101110001111110110100110100000111010101110111011100010111000001110101010101110001011100010111000101110001011100010111000111111101010111110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111011100001111111110000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111011111111111111111001111100011111000011100010111000101110001011100010111000101110001011100010111000101111001111111011000111100000111000001110101011001110001011100010111000101110001011100010111000101110001111110011111111100010111011101110111011101110111011101010111000101110001011100010111000101110001011100011111100101011101011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001010101111111111111111100111110001111100011111000111110000111000101110001011100010111000101110001011100010111000101110001010101110000011100000111000001110000011101010110011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_1 = 196'b0011110011111101111000111110111111011111000101100111111111111111111111111111111111111111111111111100011100000000000100000000000000000000100000000001111111001000000110000101000001010000000000001000;

    // Image 2: label=5, active outputs=113/196
    logic [13:0][13:0][7:0] PIXELS_2   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001111110001111100011111000111110000111100101110001011100010111000101110001011100010111000111111000111111011111111110000111000001110000011110000111111111110111000101110001011100010111000101110001011110011111111101010111011101110111010101110001011100010111000101010111111101010111000101110001011100011111100101011101011101110111010101110001011100010111000101110001011110010111100101010101011100010111000101110001010010110111010001110001011100010111000101110001011100011111100111111001111111000111000101110001011100010111000101010111111111111111100001111001011110011111100011111001111111111000011101110100011100010111000101110001011100010111000101010111100001111000011110000111100001110001011101110111011100110101110111110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111011010111010111010101110001011100010111000101110001011100010111000101111001111110011111100011111101111111011111111100000111011101010111000101110001011100010111000101110001011101011001111110000111000001110101011101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_2 = 196'b0111100111111011111111111110111111101111110111110111111111111111111111111111111111111111111111111100000000000000100000011000000001100000000000000001111111001101000001000101100000111000001000000000;

    // Image 3: label=0, active outputs=107/196
    logic [13:0][13:0][7:0] PIXELS_3   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110011111100011111000111110001111100011111000011100010111000101110001011100010111000101110001011110011111100111111101100001110000011100000111000001110111011011110001011100010111000101110001011100010111100111111101100101110111011101110101011100010111000101111011000111110111010101110001011100010111000111111001011110010101011101110101011100010111000101110001011100011111100101010101011101010111000101110001011100011111100100011101011101010111000101110001011100010111000111111001010111010101011001110001011100010111000101110001010101110101010001110001011100010111000101110001111110011111110101010111011101010111000101110001011100010111000101111101011101010111000101110001111110011111100101111111010101110111010101110001011100010111000101110001111110111111111111111100111110001111110011111101111111011101011101110101011100010111000101110001011100010111000101110001000001111111110011111111000001110000011101110111011101010111000101110001011100010111000101110001011100010111000101010101000001110101011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_3 = 196'b0011110011111111111111111111111111111111100011000111111111111111111111111111111111111111111110111100000000000000000000000000001100000000000000000001111111001100100000010001110011110000000000000000;

    // Image 4: label=0, active outputs=97/196
    logic [13:0][13:0][7:0] PIXELS_4   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110001111110111111100111100010111000101110001011100010111000101110001011100010111000101110001111110011111100110001111100001111100111111111000011100010111000101110001011100010111000101110001011100010111000111111001110011110000011100010111000101110101011111110101011100010111000101110001011100010111000101110001111110011100111100010101011101110111000101110011000111010111010101110001011100010111000101110001011100010111000111111001100011010101011001110001011100010111001100011101011101010111000101110001011100010111000101110001111110111100110100010100011101010111000101110001011100110001110101110101011100010111000101110001011100010111000101110011000011110111010101110001011100010111000101110011000111010111010101110001011100010111000101110001011100010111000111011111111111000111000101110001011100011111100101011101011101010111000101110001011100010111000101110001011100010111001110001111111111001111100011111100111111110101010001110101011100010111000101110001011100010111000101110001011100010101011100000111000001110000011101010111010101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_4 = 196'b0011100011111001111101111110111111001111100111100111111111111111111111111111111111111111111111111100000000000000000000000000000000000000010000000001111111001010000000000100000001110000000000000000;

    // Image 5: label=1, active outputs=85/196
    logic [13:0][13:0][7:0] PIXELS_5   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111001111111000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011100110101010100011100010111000101110001011100010111000101110001011100010111000101110001011100011111100101111101000001110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010100110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111101111001101000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010100110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111001101000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111111110001010101110111011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111011110101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010001111101110111011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_5 = 196'b0001100001111000111100111100011110001110000111000111111111111111111111111111111111111111111101111100001000000000000000000000000010000001000000000001111111000000000010000001000001000000000000000000;

    // Image 6: label=8, active outputs=89/196
    logic [13:0][13:0][7:0] PIXELS_6   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011110010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110011111111111111100011100010111000101110001011100010111000101110001011100010111000101110001011100011111100110011111000011110101010001110001011100010111000101110001011100010111000101110001011100010111000111111001010111010111011101010111010101000111000101110001011100010111000101110001011100010111000101110001011100010100101101010100111110011111110101110101011100010111000101110001011100010111000101110001011100010111000101110001010101111111011111111100111111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011111110001111111010111111100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010101111101111111110101011100010111000101110001011100010111000101110001011100010111000101110001111110011101110101110101011110110111110101110001011100010111000101110001011100010111000101110001011100010111000111111101010101101111100101111101110101110111000101110001011100010111000101110001011100010111000101110001011100010111000101111111111111110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_6 = 196'b0011000011110001111000111100011110001111000011100111111111111111111111111111111111111111111110111100011000000000001000000000000000000000000000000001111111000000000011000010000001010000010000000000;

    // Image 7: label=4, active outputs=94/196
    logic [13:0][13:0][7:0] PIXELS_7   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001111111000111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111110011000110101010110011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111001101010101110111010101110001011100010111000101110001011100010111000101110001111111011111110111111000111110010111010101111101011100010111000101110001011100010111000101110001011100010111000101110001010101110000011100000111110011111111111011110100011100010111000101110001011100010111000101110001011100010111000101111011010011010101011101110111000001110101011001110001011100010111000101110001011100010111000101110001011100011111100100000111011101011111100100010101011101010111000101110001011100010111000101110001011100010111000111111001010111010111010101110101000101010111011101110001011100010111000101110001011100010111000101110001111110011111110100010101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101111101000111110111011101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_7 = 196'b0001100001111001111100111110111111011111001110000111111111111111111111111111111111111111111011111100001000000000011000000000000000000000000000000001111111000100001101000000000001000001000000000000;

    // Image 8: label=3, active outputs=106/196
    logic [13:0][13:0][7:0] PIXELS_8   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111000111110001111000101110001011100010111000101110001011100010111000101110001011100010111100111111000111111111000111100010110011101010111000101110001011100010111000101110001011100010111000111111001111110011000111100000111000001110001011101110101011100010111000101110001011100010111000101110001011100010111001100001111010001100111111101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010001011110001111111111101111110011111001011100010111000101110001011100010111000101110001011100010111000101110001011101110111111100000110100011101111111011110101011100010111000101110001011100010111000101110001011100010111000111111001110011110000011100000111000001110111010101110001011100010111000101110001011100010111000101110001111110011111111100000111000101111111111111111100011110010111000101110001011100010111000101110001011100010111000101011111000001111111110011111000111110001111111111111100011100010111000101110001011100010111000101110001011100010111011100000111000001110000011000000111000001110101011001110001011100010111000101110001011100010111000101110001011100010111011100010111000001110001011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_8 = 196'b0111100011111001111100111110011111001111100111110111111111111111111111111111111111111111111111111100111000001000000000000011000000000001010000000001111111001000000011000010000001110000100000000000;

    // Image 9: label=4, active outputs=100/196
    logic [13:0][13:0][7:0] PIXELS_9   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011110010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111100111111100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010011010101011001110001011100010111000101110001011100010111000101110001011100010111000101110001111110010101110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001011101010111110101111001011110010111100101110001011100010111000101110001011100010111010111111101111110011000111111001111111111111111111011111110111111001111000101110001011100010111000101110001011100010111111100000111010101110111011101110111000011110000011100000111011101010111000101110001011100010111000111111011010011010101011001110001011100011111100110001101010101110111010101110001011100010111000101110001011100010111000101010111011101010111000101111001110111110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001111110011111110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101011111000101010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_9 = 196'b0011100001110011111101111111111111101111100011100111111111111111111111111111111111111111111111111100011000000000000010000000000000000000000000000001111111000000001011100000000001110000000000000000;

    // Image 10: label=0, active outputs=95/196
    logic [13:0][13:0][7:0] PIXELS_10   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110011111111011111000011100010111000101110001011100010111000101110001011100010111000101110001011110011111100110001101000001110101011111110101011100010111000101110001011100010111000101110001011100010111000111111001100011010101011101110111000111010111010101110001011100010111000101110001011100010111000101110001111110111100110100010100011101010111001100011101011101010111000101110001011100010111000101110001011100010111000101110011000111010111010101110001011100110001110101110101011100010111000101110001011100010111000101110001011100010111001100011101011101010111000101111011010111010111010101110001011100010111000101110001011100010111000101110001011100110101110101110101011100011111101110011111011101010111000101110001011100010111000101110001011100010111000101110011100011111111010001110001010010110001011101110101011100010111000101110001011100010111000101110001011100010111000100010111111111111111100001011111000101010111010101110001011100010111000101110001011100010111000101110001011100010111011100010111010101110111010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_10 = 196'b0011000011111001111100111110011111001111100111100111111111111111111111111111111111111111111111111100010000000000000000000000000000000000000000000001111111000010000110000001100001000000010000000000;

    // Image 11: label=7, active outputs=110/196
    logic [13:0][13:0][7:0] PIXELS_11   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110001111100001110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101010101100111000101110001011100010111000101110001011100010111000101110001011110011111100111111000111111111111111011111100111111000111000101110001011100010111000101111001111110001111100011111001111111101000111100000111100011110000011101110111011100010111000101110001011100010101010100000111000001110000011100000111010101110111011101110111011101010111000101110001011100010111000101110001011100010111000101111001111111010001010001110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111110100000111011101110111000101110001011100010111000101110001011100010111000101110001011100010111000111111000011100010111010101110001011100010111100101111001011110010111100101111001011100010111000101110001111111011111110111110111111111011111110111111101111111111111111011111110111111111111110001110001011100010111000101110111010101110111000101110111011101110001011100010111000001110000011100010111011101110111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_11 = 196'b0001110111111011111101111110111111111111110001100111111111111111111111111111111111110111111111111100001000000000000000000000001111110000000000000001111111001111000000000010000111111000000000000000;

    // Image 12: label=0, active outputs=108/196
    logic [13:0][13:0][7:0] PIXELS_12   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101111001011110010111100101111001011100010111000101110001011100010111000101110001011100010111000111111001111110011111111011111110111111101111110011110001011100010111000101110001011100010111000101111001111110011111111110001111000001110000011100000111110011101111010001110001011100010111000101110001111110011111100111001111000001110101011101110111011101010100111100000110010101000111000101110001011100011111100111111001110011110000011101110111011101010111000101110001010010110000011101010100011100010111000101110001111110011100111100010101011101110111000101110001011100010111100111111001000101100111010101110001011100010111000101001011000001110111010001110001011100010111000101111001111110011000111100000111011101010111000101110001011100010101011110001111111101000111100101111001111110011111100111001111000001110111010101110001011100010111000101110001011100010000011111001111111111101111111011111110100011110000011101010111011101010111000101110001011100010111000101110001011100010101011100000111000001110000011100000111010101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110111010101110111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_12 = 196'b0011110111111111111011111111111111101111100011100111111111111111111111111111111111111111111110111100011100000000100000000100000000000000100000000001111111011000001001000000100011100000000000000000;

    // Image 13: label=3, active outputs=103/196
    logic [13:0][13:0][7:0] PIXELS_13   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110010111100101111001011110010111100101110001011100010111000101110001011100010111000101110001011110011111100111111101111111111111111111111110111111001111100011111000011100010111000101110001011100010111000111111011100111110001011101010111000101110000011100000111000001111001010101110101011100010111000101110001011100010100101101010100011100010111000101110001011100010111000101110111010101010111000101110001011100010111000101110001010111110111010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110011111111111111010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111111111011111100001111001011110010111000101110001011100010111000101110001011100010111000101110001011100011111100111111011110011111111111111111100011100010111000101110001011100010111000101110001011100010111000111111001111111011000011100010111011101110111011001110001011100010111000101110001011100010111000101110001011100010100101111111100111110001111100011111001111111000111000101110001011100010111000101110001011100010111000101110001010101110000011100000111000001110000011101010110011100010111000101110001011100010111000101110001011100010111000101110001011101110111011101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_13 = 196'b0111110011111101111110111000011110001111000111100111111111111111111111111111111111111111111111111100111000000000001000000000000000000001100000000001111111000000101100000011100000010000000000011000;

    // Image 14: label=3, active outputs=120/196
    logic [13:0][13:0][7:0] PIXELS_14   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101111001011100010111100101111001011110010111000101110001011100010111000101110001011110011111100011111000111111111111110011111000111111111111111111111101011101010111000101110001011100010111100111111001110011110000011100000111000001110000011100000111000101110111011101110101011100010111000111111001111110011000111100010111011101110111010101110101011101010111000101110001011100010111000101110001011100010111000100000111110011111111110011111000111110001111100101111001011110010111000101110001011100010111000101110001011100010111011100010111000001110000011110001110111111101111111011111101111101010111000101110001011100010111000101110001011100010111000101111111010011110000011100000111000001110101011101110101011100010111000101110001011100010111000101110001111110011111111110001101010101110111010101110001011100010111000101110001011100010111000101110001011100010111000111111111100011111111110011111000011110010111000101110101111111010111000101110001011100010111000101110001011100010111011100000111000001111100111111111100111110001111100011111101111111001111000101110001011100010111000101110001011100010111000101110111000101110000011100000111000001110000011100000111011101010111000101110001011100010111000101110001011100010111000101110001011100010111011101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_14 = 196'b0111110111111111111111111110011111001111110011111111111111111111111111111111111111111111111110111100011101001000000000000000000000000000011000000001111111011001100111100010010001101100000010000110;

    // Image 15: label=5, active outputs=99/196
    logic [13:0][13:0][7:0] PIXELS_15   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001111110001111100101110001011100010111000101110001011100010111000101110001011100011111100111111001111111111001111100000111111111110111010001110001011100010111000101110001011100010111000111111001111111011001011101110111011101010111000101110001011101010111000101110001011100010111000101110001111110110100110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001000001111111110011111000111110001111100001110001011100010111000101110001011100010111000101110001011100010111000101110111000101110000011100000111000011111101010001110001011100010111000101110001011100010111000101110001011100010111100101111001111110011111110100000111011101010111000101110001011100010111000101110001011110011111110011111101110111111000011110001111100101110111011101110001011100010111000101110001011100010111000101010101000101110111011101110101011100010111010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_15 = 196'b0001110011111001111110111100111111011111000000000111111111111111111111111111111111111111111111111100000000001000000000001010000110000000000000000001111111001111000000000010000011110000000000000000;

    // Image 16: label=3, active outputs=113/196
    logic [13:0][13:0][7:0] PIXELS_16   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100111111000111110001111100011111000011110010111000101110001011100010111000101110001011100010111000111111001111110011000111100000111000001111100111111111111111100010111000101110001011100010111000101110001011100010111001100001101010101110111011101110111011101110001011101010101011100010111000101110001011100010111000101110001011100110100111111110100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001000101111111111011111000011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111000001111111111111111100111110001111110011110101011100010111000101110001011100010111000101110001011100010111000101110001011111110000011100000111000101110111010101110001011100010111000101110001011100010111000101110001011100011111100111111101000101110111011101110001011100010111000101110001011100010111000101110001011100010111000101110001010010110111010101111101011110010111100101111001111110001111100011110001011100010111000101110001011100010111000101011111110011111111111011111110111111111111111111001111000101110111010101110001011100010111000101110001011100010111000101010111000001110000011100010111011101110111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_16 = 196'b1111100111111011111000111110011111101111110010111111111111111111111111111111111111111111111111101101111000000000000100000100000001100000000000000001111111000010000111000001100001111100001100000000;

    // Image 17: label=4, active outputs=97/196
    logic [13:0][13:0][7:0] PIXELS_17   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111110011111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100101011101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010011010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011110011111110100000111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001110011110111110001111001011110010111000101110001011100010111000101110001011100010111000101110001111110011111111110001111111111111111111111111110111101000111000101110001011100010111000101110001011100010111100111111001010101110111011111111011000011010001011101110111011100010111000101110001011100010111000101110001111110010000011101110101111110011111110101010111011101010111000101110001011100010111000101110001011100011111100111111101011101011111100101001111010101110111010101110001011100010111000101110001011100010111000111111001010111010101011101110101011100010111010101110101011100010111000101110001011100010111000101110001011100010101010101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_17 = 196'b0001100001111001111000111110111111011111001110000111111111111111111111111111111111111111111111111100011000000000000110000000001000000000000000000001111111000000000011100010110010000000000000000000;

    // Image 18: label=6, active outputs=95/196
    logic [13:0][13:0][7:0] PIXELS_18   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111000111110000111100101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111111111001111111111111111010001110001011100010111000101110001011100010111000101110001011100011111100111001111000001110101011100010111011101110111000101110001011100010111000101110001011100010111000101110001111110110000011100000111111101000111000101001111111101000111000101110001011100010111000101110001011100010111000101001011111111001111110101010100011100010100111111110100011100010111000101110001011100010111000101110001011100010101011100000111000001110111010101110001010010110101010001110001011100010111000101110001011100010111000101110001011100010101011101110111011101010111000101001011010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111100101010100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001110011110101010001110001011100010111000101110001011100010111000101110001011100010111000101110001111111011111111100000111011101110111000101110001011100010111000101110001011100010111000101110001011100010111000101110111000101110111011101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_18 = 196'b0011000011110001111000111110011110000111100011110111111111111111111111111111111111111111111111111100000000011000000000000100000000000000000000000001111111001110000100000010000000110000011000000000;

    // Image 19: label=1, active outputs=85/196
    logic [13:0][13:0][7:0] PIXELS_19   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111011111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110100000111011101010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001000001110111010101110001011100010111000101110001011100010111000101110001011100010111000111111001111110011000111101010111011101010111000101110001011100010111000101110001011100010111000101110001011100011111100111001111000101010111010101110001011100010111000101110001011100010111000101110001011100010111000111111001110011110000011101010110011100010111000101110001011100010111000101110001011100010111000101110001011100011111100110001111010101110111010101110001011100010111000101110001011100010111000101110001011100010111000111111011110011110001010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111001100001101010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100110001110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011101010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_19 = 196'b0001100001111000111100111110011110001110000111000111111111111111111111111111111111111111111111111100001000000000000000000000000000000000000000000001111111000010000000000010000000000000100000000000;

    // Image 20: label=3, active outputs=107/196
    logic [13:0][13:0][7:0] PIXELS_20   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110001111100011111001011110010111000101110001011100010111000101110001011100010111000101110001011110011111110110001111100011111111111111111110111110000111000101110001011100010111000101110001011100011111100111111001000101010111011101110111011101110001011111111111111111000111010101110001011100010111000101110001011100110000111111111100111100010111000101110001011100010001011100010101011101010111000101110001011100010111000101110001000101111100111111110100011100010111000101110001011100010111010101110001011100010111000101110001011100010111000101110011000001111111111011111000011110010111100101110001011100010111000101110001011100010111000101110001011100010111000101110111010011111100111011111110111111000111000101110001011100010111000101110001011100010111000101110001011100011111100111111101000001110000011101010101011100010111000101110001011100010111000101110001011100010111000111111011110011110100011001111111011111010111100111111000011100010111000101110001011100010111000101110001011100010111000100000111100011111111111111111110111111111101111111010110011100010111000101110001011100010111000101110001011100010111011101010111000101110000011100010111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_20 = 196'b0111100111111011111110111110011110001111100110110111111111111111111111111111111111111111111111101100111000000010000000000000000001100000000000000001111111000011000010000001100001111000001100000000;

    // Image 21: label=9, active outputs=90/196
    logic [13:0][13:0][7:0] PIXELS_21   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111100111111000111100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111010000011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100100011101011101110111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010111010101011001110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110100010101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010111110111111001111001011100010111000101110001011100010111000101110001011100010111000101110001011110011111100111111100111111111111110011111000011100010111000101110001011100010111000101110001011100010111000111111011100011110000011100000111000001110101010001110001011100010111000101110001011100010111000101110001111110010111010101000111111111101111100100011111011101110111000101110001011100010111000101110001011100010111000101001111111111001111110111111111000001110111011101110001011100010111000101110001011100010111000101110001011100010101010100000111010101110111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_21 = 196'b0001110001111001111000111110011111001111000000000111111111111111111111111111111111111111111111111100011000000000000010000010000000000000000000000001111111000000000011000000000001110000000000000000;

    // Image 22: label=7, active outputs=99/196
    logic [13:0][13:0][7:0] PIXELS_22   = 1568'b01110001011100010111000101110001011100010111000111111000111110001111100001110001011100010111000101110001011100010111000101110001011100010111000101110001111110110100110110000111110111101111010101110001011100010111000101110001011100010111000101110001011100010111000101110001010101111100101100010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001010011010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001111110011100110100010100011101010111000101110001011100010111000101110001011100010111000101110001011100010111100111111101000001110111011101110001011100010111000101110001011100010111000101110001011100010111000111111001111110011000110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111101101001111000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110110111010101111110011110010111100101111001011110010111100101111001011100010111000101110001011100010111000101001011110011101111111011111111111111111111111111111111111111111111110101110001011100010111000101110001011100010101010100000111000001110001011101110111011101110111011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_22 = 196'b0011110001111001111100111110011111100111110000000111111111111111111111111111111111111111111111111100101100000000000000000010000001110000000000000001111111000000000110000010000001111000000000000000;

    // Image 23: label=1, active outputs=84/196
    logic [13:0][13:0][7:0] PIXELS_23   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110011111100001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001110111011111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111100111111001000101010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011000110101010110011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111001101000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010001010101110111011100010111000101110001011100010111000101110001011100010111000101110001011100011111100101001101011101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011000110111010110011100010111000101110001011100010111000101110001011100010111000101110001011100011111101111001101000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010001011101110111011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_23 = 196'b0001110001111000111100111100011110001110000011000111111111111111111111111111111111111111111110111100001000000000000000000000000000000000000000000001111111000011000000000001000000000000100000000000;

    // Image 24: label=5, active outputs=116/196
    logic [13:0][13:0][7:0] PIXELS_24   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111000111110001111110011111100111110001111100101110001011100010111000101110001011100010111000101111001111110001111111100000111000101110001011100000111111111111111100001110001011100010111000101110001111110011111100110001101010101110111010101110001011100010111011100000111110111111111010101110001011100010111000111111001010011010101011101110101011100010111000101110001011100010111011101010111011101010111000101110001111110011111100101010100011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001000001111111110011111000011110010111100101111001111110011111100011111000111110000111000101110001011100010111000101010111000001111100111111111110111111101111111011111110100011110000011001010100011100010111000101110001011100010111000101110111010101110000011100000111000001110000011100000111000001110101010001110001011100010111000101110001011100010111000101110001011100011111101111111000111110001111100011111001011101000111000101110001011100010111000101110001011100010111000101110001010111110000011100000111000001110000011111011111111101010111000101110001011100010111000101110001011100010111000101110111000101110001011101110111011101110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_24 = 196'b1111100111111111111111111110111111000111110011111111111111111111111111111111111111111111111110111100111101000000000000010100000000110000000000000001111111011001000000000111000001111000000100000000;

    // Image 25: label=2, active outputs=106/196
    logic [13:0][13:0][7:0] PIXELS_25   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111110010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111111011100010111000101110001011110011111100011111000111110001111100001110001011100010111000101110001011100011101111111111101111110011111100011111001100011110000011100000111110111011111010101110001011100010111000101110001011100011100011111111111110011110000011011001110111110001100111100010100011101010111000101110001011100010111000101111001111110010000011100000111000001110000011100000111000101110111011101110001011100010111000101110001011100011111101110001101010101100111000101110001011101110111010101110001011100010111000101110001011100010111000101110001010011110001010001110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101001111111101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010101111111111110111110010111100101111001011100010111000101110001011100010111000101110001011100010111000101110001011100111000111111111111111111101111110001110001011100010111000101110001011100010111000101110001011100010111000101110001011101110001011100000111010101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_25 = 196'b1100000111111101111110111111011111001111000111100111111111111111111111111111111111111111111110111100000000010001000000000001000110000000000000000001111111011001100100110000100011000000110000000000;

    // Image 26: label=9, active outputs=104/196
    logic [13:0][13:0][7:0] PIXELS_26   = 1568'b01110001011100010111000111111001111110000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010111110101010100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110011000111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111011101011101010111000101110001011110010111100101110001011100010111000101110001011100010111000101110001010010110001010101110101111110001111100111111111111111111111110001110001011100010111000101110001011100010111000101010111011111011111100101001101000101110111011101110111100101111111110101110001011100010111000101110001011100010111001100011101110011110001010101110101011100010111000101110001000001111111010001110001011100010111000101110001011100010000111111011011011111000111000101110001011100011111100111111001010101000111000101110001011100010111000101110001010101111000111111111110111110000111100111111001111110011000111101010100011100010111000101110001011100010111000101110001010101110000011111001111111111111111111110001111000001110111010101110001011100010111000101110001011100010111000101110001011100010111011100010111000101110111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_26 = 196'b1110000111110011111101111111011111001111110000000111111111111111111111111111111111111111111111111111000000001100000000000010000001000000000000000001111111000110000001100011110000110000000000000000;

    // Image 27: label=1, active outputs=88/196
    logic [13:0][13:0][7:0] PIXELS_27   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111011111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011100110100000111011101010111000101110001011100010111000101110001011100010111000101110001011100011111100111111001100011010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010100110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101000101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011110110001010101110111011100010111000101110001011100010111000101110001011100010111000101110001011100011111100101011101010101100111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010001010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011111010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_27 = 196'b0001100001111000111100111110011110011110001111000111111111111111111111111111111111111111111111111100001000000000000000000000000010000000000000000001111111000000000000000001000001000000100000000000;

    // Image 28: label=3, active outputs=97/196
    logic [13:0][13:0][7:0] PIXELS_28   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110011111100011111000011100010111000101110001011100010111000101110001011100010111000111111001111110001111110111111111100001110101010101110001011100010111000101110001011100010111000101110001111110011111110110000111010101110111011101110101011100010111000101110001011100010111000101110001011100010111000101011111011101000111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111011101000111111111000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111011110010111111111111111100001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111111010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110101010110011100010111000101110001011100010111000101110001011100010111000101110001011110011111100111011111010101110111010101110001011100010111000101110001011100010111000101110001011100010111000111111111100011111111110011111100111111000111000101110001011100010111000101110001011100010111000101110001011100010111011100010111000001110001011101110111011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_28 = 196'b0011110011111001111100111100011110001111000111100111111111111111111111111111111111111111111111111100011100000000000100000000000000000000000000000001111111001010000011000000100001100000000000000000;

    // Image 29: label=3, active outputs=101/196
    logic [13:0][13:0][7:0] PIXELS_29   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001011110010111100101111001011100010111000101110001011100010111000101110001011100010111000101111001111110011111111111111111111111111111111111110100011100010111000101110001011100010111000101110001011110010111110110010111011101110111011101110111010101110101010101110001011100010111000101110001011100011111100101111001010101110111010101110001011100010111000101110001010101010111000101110001011100010111000101110001011100110101010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001110111111111000101110001011110010111100101110001011100010111000101110001011100010111000101110001011100010111000111011111111111011111100011111111111111101111010001110001011100010111000101110001011100010111000101110001011100011111100100011111000001110000011100010111011101110111000101110001011100010111000101110001011100010111000111111001011111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010101111101110100011110010111100101111001011100010111000101110001011100010111000101110001011100010111000101110001011101111000111111111111110111111001011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_29 = 196'b0011110011111101111100111100011111001111000111100111111111111111111111111111111111111111111101111100011100000000000000000011000000000000000000000001111111000111000000000011100000100000110000000000;

    // Image 30: label=8, active outputs=92/196
    logic [13:0][13:0][7:0] PIXELS_30   = 1568'b01110001011100010111000101110001011100010111100101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111111111110011111000011100010111000101110001011100010111000101110001011100010111000101110001111110011111111110000111000001110111110011110001011100010111000101110001011100010111000101110001011100010111000101110001011111110111010111111001100111010111010101110001011100010111000101110001011100010111000101110001011100011111100111111111111110001100110100010100011101010111000101110001011100010111000101110001011100010111000101110001011100010001011110001111100011010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110111000111111111100011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111001000001110000011111111110111110000111000101110001011100010111000101110001011100010111000101110001011100110000110101110100011101110001011111111111011101000111000101110001011100010111000101110001011100010111000101110001000001111111111111111100111110001111101011011101111101010111000101110001011100010111000101110001011100010111000101110001010101110000011100000111000001110000011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_30 = 196'b0111100011110001111000111100011111000111100001110111111111111111111111111111111111111111111111111101110000000000000000000000000000000000000000000001111111001000000000000001100000110000000000000000;

    // Image 31: label=9, active outputs=100/196
    logic [13:0][13:0][7:0] PIXELS_31   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111011111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011100110100000111011101010111000101110001011100010111000101110001011100010111000101110001011100010111100111111101000001110111011101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010001010101110111011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101011111001111100011111000111110001111000101110001011100010111000101110001011100010111000101111001111110011000111011111111110011110000011100010111011101010111000101110001011100010111000101110001011100011111100110001111000001110101011101110111011111001111110101110101011100010111000101110001011100010111000101110101100011110101011101110101011110011111100011111101000101010111010101110001011100010111000101110001011100011111100111111001111110001111100011111101110011110101011101110101011100010111000101110001011100010111000101110001011100010000011110001111000001110001011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_31 = 196'b0011110001111001111101111110111111011111100111000111111111111111111111111111111111111111111111111100011100000000000000000000000000000000000000000001111111000100000110000001100001100000000000000000;

    // Image 32: label=6, active outputs=90/196
    logic [13:0][13:0][7:0] PIXELS_32   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110011111100001110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100011111001100011111111010001110001011100010111000101110001011100010111000101110001011100010111000111111001111111010000011101000111010111111111010101110001011100010111000101110001011100010111000101110001011100010111101100010101010101111111111110011111011101010111000101110001011100010111000101110001011100010111000111111011010011010101010001111011111110110001011001110101011100010111000101110001011100010111000101110001011100010111001111001101111111001111100110001111000101100111010101110001011100010111000101110001011100010111000101110001011100010000011100000111000001100000011000010101011101010111000101110001011100010111000101110001011100010111000101110001011101110001011100000111000001110101010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010100101100010101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010011110101010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101010101011101110111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_32 = 196'b0011000011110001111100111110011011001111000011100111111111111111111111111111111110111111111111111100000000000000000000000000000000000000000000000001111111000110000111000010000001000000010000000000;

    // Image 33: label=2, active outputs=115/196
    logic [13:0][13:0][7:0] PIXELS_33   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111111111111110001110001011100010111000101111001011110010111100101111001011110010111000101110001011100010111000101001111111101000111000111111001111110001111100111111110111111101111111111111100011100010111000101110001011100010100101111111100111110001111111110001111000001110000011100000110000101100111010101110001011100010111000101110001010010111000111010001111010001110111111111111111000011110000011100010111011101010111000101110001011100011111100111111001000001110000011111001111111111110101011101110111011101110111010101110001011100010111000101110001111110011100110101010111011101110111011101110111011101010111000101110001011100010111000101110001011100010111000101011111010101110111010101110001011100010111000101111001011110010111000101110001011100010111000101110001011100010111011100000111111111001111100011111000111110001111111111111100011101010111000101110001011100010111000101110001011100010101011100000111100011111000111100000111000001110001010101110101011100010111000101110001011100010111000101110001011100010111011101110111011101110111011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_33 = 196'b0101110011111111111111111111111111011111100111110111111111111111111111111111111111111111111110011101100000000010000011000100000000000000010000000001111111001111100011100110000000010000011000000000;

    // Image 34: label=8, active outputs=107/196
    logic [13:0][13:0][7:0] PIXELS_34   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110001111100011111000011100010111000101110001011100010111000101110001011100010111000101110001111110011111111111001111000001111101111111110001011100010111000101110001011100010111000101110001011100010111000111011111000001110111011001110111000001111111010001110001011100010111000101110001011100010111000101110001011100010111000100000111111111111111100001111011110111101111010101110001011100010111000101110001011100010111000101110001011100010111011100000111110011111100111100010110011101010111000101110001011100010111000101110001011100010111000101110001011110011111101110001111000001101100111011111100111100010111000101110001011100010111000101110001011100011111100011111001110011110000011100000111000001111100111111111000011100010111000101110001011100010111000111111001111111110000011000000111010101010111000101111011010011111101111011110101011100010111000101110001011101011000111100000111000001100111011011111101111110001111100110001111000101110111010101110001011100010111000101110001011101110000011100000111110011111111111110001111000001110001011101110101011100010111000101110001011100010111000101110001011100010111011101010111011101110111011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_34 = 196'b0111000011110001111101111110111111111111110111110111111111111111111111111111111111111111111111011100110000001000011000000000000110000000000000000001111111001100000000000100010000110001010000000000;

    // Image 35: label=7, active outputs=109/196
    logic [13:0][13:0][7:0] PIXELS_35   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110111110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101010101110111010101110001011100010111000101110001011100010111000101110001011100010111000111111001010111010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001111110011111100111111100111110001111100011111000011100010111000101110001011100010111000101111001111110001111100011111101100011110000011100000111000001110101010101110001011100010111000101110001011100010101010100000111000001110000011101110111011101110111011101110101011100010111000101110001011100010111000101110001111110011111100100011111011101110111000101110001011100010111000101110001011100010111000101110001011100010111000111111001000111010111011101110001011100010111100111111001111110000111000101110001011100010111000101110001111110110100110101110100011110010111100111111001111110011111111011011101111101010111000101110001011100010111000101110011100001111111011111111111111111111100111100000111000001110101011101110101011100010111000101110001011100010111000101110101011101010111011101110111011100010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_35 = 196'b0001110001111011111101111100111111011111101111100111111111111111111111111111111111111111111101111100011100000000000110001000001010000000000000000001111111000100000000000110100011111000110000000000;

    // Image 36: label=9, active outputs=86/196
    logic [13:0][13:0][7:0] PIXELS_36   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010010110101010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111111010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110110101110101110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111001110111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111111010100111110000111011101111111000101110001011100010111000101110001011100010111000101110001011100010111000101110111000101110111011101001111111101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110010111110101010100011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111111001000111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100111100111100010101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_36 = 196'b0011100001110001111000111100011110000111000011100111111111111111111111111111111111111111111111111100111000000000000000000000000000000000000000000001111111000100000110000000000000000000000000000000;

    // Image 37: label=7, active outputs=107/196
    logic [13:0][13:0][7:0] PIXELS_37   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110111110101011100010111000101110001011100010111000101110001011100010111000101110001011100011111100111001101000001110111010101110001011100010111000101110001011100010111000101110001011100010111000101111001111110010111010111111110011100010111000101110001011100010111000101110001011100010111100101111001111110001111100110001111110011101100111111110100011100010111000101110001011100010111000111111101111111111111111111001111000001110000011100000111000101110111011101110001011100010111000101110001011100010111000101110111111110110000110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101010101110111010101110001011100010111000111111001111110000111000101110001011100010111000111111001011111010001010001110101011100010111100111111001111110001111111101010100011100010111000101110001011100011111100111001101111111001111100011111000111111011111111110001111000001110101010101110001011100010111000101110001010111110000011100000111000001110000011100010111011101110111011101110101011100010111000101110001011100010111000101110001011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_37 = 196'b0001110011111011111101111111111111011011100110000111111111111111111111111111111111111111111101111100011100000000011000000000000000010001000000000001111111000011001100000001110010110000100000000000;

    // Image 38: label=9, active outputs=103/196
    logic [13:0][13:0][7:0] PIXELS_38   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111101111111001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100110101110111110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110011000111010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111001111001101111111011111110111111101111111011111100001110001011100010111000101110001011100010111000101110001011100110000110101010111011101110111011101110111010001111111110011110001011100010111000101110001011100010111000101111011010101010111010101110001011100010111000101110111000011111111010001110001011100010111000101110001011100011111101101010100011100010111000101110001011100010111000101110111010101000111000101110001011100010111000101110001010010110101010001110001111111111111010101110001011100011111111101010100011100010111000101110001011100010111000101011111010101010111000111111111111111000111100111111000111111010111010101110001011100010111000101110001011100010111000101110101011100010111011110001111111111111001111101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_38 = 196'b0110000011110001111100111111011111001111110001110111111111111111111111111111111111111111111111111101100000011100000000000010000100000000000000000001111111001110000011000001000000111000000000000000;

    // Image 39: label=9, active outputs=98/196
    logic [13:0][13:0][7:0] PIXELS_39   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111111011111010001110001011100010111000101110001011100010111000111111101111111010111000101110001011100011111100100011101011101110111000101110001011100010111000101110001011100010111100101111101011100010111000111111001111111010101011001110001011100010111000101110001011100010111000101110001110111011101010101110001111110010111100101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001000111110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111100111111100111110001111100001110001011100010111000101110001011100010111000101110001011100010111000101111011110011011101111110000111000001111111010001110001011100010111000101110001011100010111000101110001011100011111100100000111011111111111100101011101011101110111000101110001011100010111000101110001011100010111000111111011110011011111110011111101100111110101010101110001011100010111000101110001011100010111000101110001011100010111001100001111000001110001011101110111011100010111000101110001011100010111000101110001011100010111000101110001011100010111011101110111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_39 = 196'b1101100111111011111000111100011111001111000111000111111111111111111111111111111111111111111111111101011000000000000000000000000010000000000000000001111111011100000000000011000001100000000000000000;

    // Image 40: label=8, active outputs=99/196
    logic [13:0][13:0][7:0] PIXELS_40   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111100011111000011110010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101100001111000011111111101111100010111000101110001011100010111000101110001011100010111000111111011010011010101011101110101011100010100111111110100011100010111000101110001011100010111000101110001011100010111001101001111111110000111000111111001010111010101011001110001011100010111000101110001011100010111000101110001011100010101011111111111111111001111110100010101011101010111000101110001011100010111000101110001011100010111000101110001011100010111111100000110100011101111110001111001011100010111000101110001011100010111000101110001011100010111000111111001110011010000011100000111100011111111111011110001011100010111000101110001011100010111000101110001011100011111100100000111011101110111000101111011010111110111010101110001011100010111000101110001011100010111000111111001010111110111010011111001111110001111110100000111011101010111000101110001011100010111000101110001011100010111000101001111111111001111110100000111000101110111011101110001011100010111000101110001011100010111000101110001011100010101010100000111010101110111011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_40 = 196'b0111100011111001111000111110011111001111100001100111111111111111111111111111111111111111111111011100111000000000000100000100000000000000000000000001111111000010000110000010110001100000010000000000;

    // Image 41: label=4, active outputs=95/196
    logic [13:0][13:0][7:0] PIXELS_41   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110001111100001110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111100101001101010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111111010000011101110101011100010111000101110001011100010111000101110001011100010111000101110001011110011111100111001111011111000111000101110001011100010111000101110001011100010111000101110001011100011111110111111001110011111000111011111110111111000111000101110001011100010111000101110001011100010111000101110001011110110100111100000111000001110000011100000111110101100111000101110001011100010111000101110001011100010111000111111001000101010111111011111000010011010101011101110101011100010111000101110001011100010111000101110001111110010100110101110100111110011000110101010111011101010111000101110001011100010111000101110001011100011111100111111101000001110101010110001111010101110111010101110001011100010111000101110001011100010111000101110001011100110000110101110101011100010111010101110101011100010111000101110001011100010111000101110001011100010111000101110001010101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_41 = 196'b0001110001110001111100111110111111011111000110000111111111111111111111111111111111111111111111111100001000000000000010000001000000000000000000000001111111000100000111000001100010000000000000000000;

    // Image 42: label=4, active outputs=102/196
    logic [13:0][13:0][7:0] PIXELS_42   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101111111011111010001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101001111010101000111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111100101110100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111011010011111101010001110101011110010111100101110001011100010111000101110001011100010111000101110001011100011111101110001111111111101111110011111001111111001111100001110001011100010111000101110001011100010111000101110001010010110000011000000111000001110000011100000111111111001111000101110001011100010111000101110001011100010111100111111001000001110001011101110111011101110000111100010110011101010111000101110001011100010111000101110001111110011000111100010100011101010111000111111001110011110001010101110101011100010111000101110001011100011111101111001111000101010111011101110001111110111100111100000111010101100111000101110001011100010111000101110001011100010001011101010101011100010111000101110011000011110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_42 = 196'b0111000011110001111100111111111111111111100001110111111111111111111111111111111111111111111111111100110000000000000000000100000000000000000000000001111111001000000111000011100001010000000000000000;

    // Image 43: label=2, active outputs=102/196
    logic [13:0][13:0][7:0] PIXELS_43   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001111110011111110001110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101011111011101000111000101110001011100010111000101111001011110010111100101111001011100010111000101110001011100010111001111111111111110000111100111111000111110011111111111111110111111111111110001110001011100010111000101110001011100010101011111001111111111111100111100000111000011110000011100010111011101110111000101110001011100010111000101111001111111010001111100010111011101110111011101110111011101110111010101110001011100010111000101110001011110010111110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000111111011010101010111010101110001011110010111100101110001011100010111000101110001011100010111000101110001011100010101011111111111111110001111100011111111110111110111010101110001011100010111000101110001011100010111000101110001011100010101011100000111000001110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_43 = 196'b0100000011111001111111111111111110011111000111000111111111111111111111111111111111111111111111111100000000000110000010000000000001000000000000000001111111001011100110010000000010110000000000000000;

    // Image 44: label=5, active outputs=105/196
    logic [13:0][13:0][7:0] PIXELS_44   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110001111100011111000111110010111000101110001011100010111000101110001011100010111000101110001111110011111100110001111000001111000111111111110111110000111000101110001011100010111000101110001011100010111100111111001000001110000011101010111010101110000011111011110111101010111000101110001011100010111000101110001111110111000111101010100011101010111000101110001011110110001011101110101011100010111000101110001011100010111000101001011000001100101010001110001011100011111100111001111000101010111010101110001011100010111000101110001011100010101011100000111011101000111100101110001011110011111101111111000011100010111000101110001011100010111000101110001011100010001011111001111111111001111100011111001111111101000111111110100011100010111000101110001011100010111000101110001011100010101011100000111000001110000011100000111000001110101010001110001011100010111000101110001011100010111000101110101111111011111100101111101111110001111100100010110011101010111000101110001011100010111000101110001011100010111000101001111111111101111111011001111000001110001011101110101011100010111000101110001011100010111000101110001011100010101010100000111000001110001011101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_44 = 196'b0111100111111011111101111110011111001111100001110111111111111111111111111111111111111111111111111100111000000000000000000000000011000000000000000001111111000011000001000110100001110000000000000000;

    // Image 45: label=5, active outputs=106/196
    logic [13:0][13:0][7:0] PIXELS_45   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110011111100011111000111110001111100001110001011100010111000101110001011100010111000101110001011110011111100111111111100011111000011100000111010101100111000101110001011100010111000101110001011100011111100111111101000001110101011101110111011100010111011101110101011100010111000101110001011100010111000101110001011100110100110101111100011110010111100101111001011110010111100101110001011100010111000101110001011100010111000101110001000001111111111111111111111111111111111111111110110111000111010101110001011100010111000101110001011100010111000101110001010101110001011101110111011111110000011101010110011100010111000101110001011100010111000101110001011100010111100111111001111110001111100011111101010101110111010101110001011100010111000101110001011100011111100011111000111111111111111110001111000001110101011101110101011100010111000101110001011100010111000111111001111111010000011101010111011101110111011101110111011101010111000101110001011100010111000101110001011101011000111101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011101010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_45 = 196'b0011100011111001111100111111111111011111101110000111111111111111111111111111111111111111111111111100000000000000000110000000001010000000000000000001111111001100000111100001100011100001000000000000;

    // Image 46: label=4, active outputs=95/196
    logic [13:0][13:0][7:0] PIXELS_46   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011110010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100011111101111111101111100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100111000111111110100011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110011000011110101010001110001011110011111100001110001011100010111000101110001011100010111000101110001011100010111101101011101111111001111100011111101100011111111110001110101011100010111000101110001011100010111000101110001111110011100011111111111100111110101011101001111000101000111010101110001011100010111000101110001011100011111100111001111100011011001011101110111011110110101110101110101011100010111000101110001011100010111000101110001111110011000110101010111011101010111000111111001000001110111010101110001011100010111000101110001011100010111010110001111010101110111010101110001111110010101110101110101011100010111000101110001011100010111000101110001011100010111010101110101011100010111000111111111000001110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011101010111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_46 = 196'b0110000011110001111100111111111111011111100001100111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000001111111001100000111100000000000010000000000000000;

    // Image 47: label=8, active outputs=104/196
    logic [13:0][13:0][7:0] PIXELS_47   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101111001111110001111100011111000111100010111000101110001011100010111000101110001011100010111000101110001011110011111110111001111000001110100011111110100011100010111000101110001011100010111000101110001011100010111000111111111000001110111011111111001010011010111010101110001011100010111000101110001011100010111000101110001111110010111110101110100111110001111110101010111011101010111000101110001011100010111000101110001011100010111000101110001010011111111110011111101010101110111010101110001011100010111000101110001011100010111000101110001011110011111100111111111000001110101011101110101011100010111000101110001011100010111000101110001011100011111100011111101100111110000011101111101111100010111000101110001011100010111000101110001011100010111000111111101111111010001011101110111011110110001110101110101011100010111000101110001011100010111000101110001011100010111011101010111011111011111100011111101000101010111010101110001011100010111000101110001011100010111000111111001111111011111100011111101100111110001011101110111011100010111000101110001011100010111000101110001011100010111000101010111000001110101011101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_47 = 196'b0011110001111101111111111110111110011111001111000111111111111111111111111111111111111111111111111100011100000000001000000000001000000000000000000001111111000111000000000111000010100000000000000000;

    // Image 48: label=9, active outputs=101/196
    logic [13:0][13:0][7:0] PIXELS_48   = 1568'b01110001011100010111000101110001011100010111100101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111011111111011111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111001100011101011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100110101010101110101011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001011111010111100101111001011110010111100101110001011100010111000101110001011100010111000101110001011100010100101111111100111111011101111111111111111111111111010001110001011100010111000101110001011100010111000111111001111110010000011101010111011101010111011101110111010101000111000101110001011100010111000101110001011100010111101100011101010101100111000101110001111110010111100111010101011100010111000101110001011100010111000101110001111110110101010101110101011100010111100111111001000111110111010101110001011100010111000101110001011100010111000101010111111111011111100111111001111111011001111101110111011100010111000101110001011100010111000101110001011100010111000100000111111111111111111101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101110111011101110111010101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_48 = 196'b0111000011110001111100111110011111001111100011100111111111111111111111111111111111111111111110111101110000000000000110000000000010000000000000000001111111000000000111100010000011110000010000000000;

    // Image 49: label=6, active outputs=92/196
    logic [13:0][13:0][7:0] PIXELS_49   = 1568'b01110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111100111111000011100010111000101110001011100010111000101110001011100010111000101110001011100010111000111111001111110011111110011111000111110000111000101110001011100010111000101110001011100010111000101111001111110001111110110001111000001110000011101010100011100010111000101110001011100010111000101110001011110011111100110001101000101110111011101111111010011010101010001110001011100010111000101110001011100011111100111111001100011010101011101110101011100011111100100010101011101010111000101110001011100010111000101110001011100110000111101010111011101010111000111111001111111010101011001110001011100010111000101110001011100010111000101110001011101010111010101110001111110011111110101010111011101010111000101110001011100010111000101110001011100010111000101110001011100011111100111111101010101110111010101110001011100010111000101110001011100010111000101110001011100010111100111111000111111010101011101110101011100010111000101110001011100010111000101110001011100010111000101110001111111110000011101010111011101010111000101110001011100010111000101110001011100010111000101110001011100010111000101010101011101110111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001;
    logic [3:0][6:0][6:0]   EXPECTED_49 = 196'b0001000011111011111101111110111111001111000111000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111000110000001000000100000000001000000000000;

    // DUT signals — multi-dimensional types matching layer_two.sv ports
    logic [13:0][13:0][7:0] pixels;
    logic [2:0][2:0][7:0]   weights;
    logic [3:0][6:0][6:0]   layer_two_out;
    logic done, clk, rst_n;
    state_t state;

    // Module-level staging regs — avoids multi-dim task params (icarus 10.2 limitation)
    logic [13:0][13:0][7:0] test_pixels;
    logic [3:0][6:0][6:0]   test_expected;

    integer errors = 0, total_checks = 0;

    layer_two dut (
        .clk(clk), .rst_n(rst_n), .state(state),
        .pixels(pixels), .weights(weights),
        .layer_two_out(layer_two_out), .done(done)
    );

    initial begin clk = 0; forever #5 clk = ~clk; end

    // ================================================================
    // run_test: drives DUT and compares using [filter][row][col] indexing
    //           — no flat bit manipulation, purely multi-dim access
    // ================================================================
    // run_test: uses module-level test_pixels/test_expected (set before each call).
    //   Comparison loop uses computed flat bit index [f*49+r*7+c] — equivalent
    //   to [f][r][c] for a [3:0][6:0][6:0] array but supported by icarus 10.2.
    //   Declarations remain multi-dim throughout.
    task run_test;
        input integer img_idx, label;
        integer f, r, c, bit_pos, mismatches;
        begin
            mismatches = 0;
            rst_n = 0; state = s_IDLE;
            pixels  = test_pixels;
            weights = TRAINED_WEIGHTS;
            #20; rst_n = 1;
            #20; state = s_LAYER_2;
            wait(done == 1);
            #100;

            // bit_pos = f*49 + r*7 + c  (same as [f][r][c] for [3:0][6:0][6:0])
            for (f = 0; f < 4; f = f + 1)
                for (r = 0; r < 7; r = r + 1)
                    for (c = 0; c < 7; c = c + 1) begin
                        bit_pos = f*49 + r*7 + c;
                        total_checks = total_checks + 1;
                        if (layer_two_out[bit_pos] !== test_expected[bit_pos]) begin
                            mismatches = mismatches + 1;
                            errors     = errors + 1;
                        end
                    end

            if (mismatches == 0)
                $display("PASS  image=%0d  label=%0d  (196/196 outputs correct)", img_idx, label);
            else
                $display("FAIL  image=%0d  label=%0d  (%0d/196 mismatches)", img_idx, label, mismatches);
        end
    endtask

    initial begin
        $dumpfile("layer_two.vcd");
        $dumpvars(0, tb_layer_two);

        $display("\n====================================================");
        $display("Layer Two vs Reference Model");
        $display("Inputs:    layer_one output on real MNIST images");
        $display("Weights:   derived from layer_3_weights.mem (majority vote)");
        $display("Threshold: 41 42 35 37 (from layer_4_thresholds.mem)");
        $display("Testing 50 images");
        $display("====================================================\n");

        test_pixels   = PIXELS_0;
        test_expected = EXPECTED_0;
        run_test(0, 5);

        test_pixels   = PIXELS_1;
        test_expected = EXPECTED_1;
        run_test(1, 3);

        test_pixels   = PIXELS_2;
        test_expected = EXPECTED_2;
        run_test(2, 5);

        test_pixels   = PIXELS_3;
        test_expected = EXPECTED_3;
        run_test(3, 0);

        test_pixels   = PIXELS_4;
        test_expected = EXPECTED_4;
        run_test(4, 0);

        test_pixels   = PIXELS_5;
        test_expected = EXPECTED_5;
        run_test(5, 1);

        test_pixels   = PIXELS_6;
        test_expected = EXPECTED_6;
        run_test(6, 8);

        test_pixels   = PIXELS_7;
        test_expected = EXPECTED_7;
        run_test(7, 4);

        test_pixels   = PIXELS_8;
        test_expected = EXPECTED_8;
        run_test(8, 3);

        test_pixels   = PIXELS_9;
        test_expected = EXPECTED_9;
        run_test(9, 4);

        test_pixels   = PIXELS_10;
        test_expected = EXPECTED_10;
        run_test(10, 0);

        test_pixels   = PIXELS_11;
        test_expected = EXPECTED_11;
        run_test(11, 7);

        test_pixels   = PIXELS_12;
        test_expected = EXPECTED_12;
        run_test(12, 0);

        test_pixels   = PIXELS_13;
        test_expected = EXPECTED_13;
        run_test(13, 3);

        test_pixels   = PIXELS_14;
        test_expected = EXPECTED_14;
        run_test(14, 3);

        test_pixels   = PIXELS_15;
        test_expected = EXPECTED_15;
        run_test(15, 5);

        test_pixels   = PIXELS_16;
        test_expected = EXPECTED_16;
        run_test(16, 3);

        test_pixels   = PIXELS_17;
        test_expected = EXPECTED_17;
        run_test(17, 4);

        test_pixels   = PIXELS_18;
        test_expected = EXPECTED_18;
        run_test(18, 6);

        test_pixels   = PIXELS_19;
        test_expected = EXPECTED_19;
        run_test(19, 1);

        test_pixels   = PIXELS_20;
        test_expected = EXPECTED_20;
        run_test(20, 3);

        test_pixels   = PIXELS_21;
        test_expected = EXPECTED_21;
        run_test(21, 9);

        test_pixels   = PIXELS_22;
        test_expected = EXPECTED_22;
        run_test(22, 7);

        test_pixels   = PIXELS_23;
        test_expected = EXPECTED_23;
        run_test(23, 1);

        test_pixels   = PIXELS_24;
        test_expected = EXPECTED_24;
        run_test(24, 5);

        test_pixels   = PIXELS_25;
        test_expected = EXPECTED_25;
        run_test(25, 2);

        test_pixels   = PIXELS_26;
        test_expected = EXPECTED_26;
        run_test(26, 9);

        test_pixels   = PIXELS_27;
        test_expected = EXPECTED_27;
        run_test(27, 1);

        test_pixels   = PIXELS_28;
        test_expected = EXPECTED_28;
        run_test(28, 3);

        test_pixels   = PIXELS_29;
        test_expected = EXPECTED_29;
        run_test(29, 3);

        test_pixels   = PIXELS_30;
        test_expected = EXPECTED_30;
        run_test(30, 8);

        test_pixels   = PIXELS_31;
        test_expected = EXPECTED_31;
        run_test(31, 9);

        test_pixels   = PIXELS_32;
        test_expected = EXPECTED_32;
        run_test(32, 6);

        test_pixels   = PIXELS_33;
        test_expected = EXPECTED_33;
        run_test(33, 2);

        test_pixels   = PIXELS_34;
        test_expected = EXPECTED_34;
        run_test(34, 8);

        test_pixels   = PIXELS_35;
        test_expected = EXPECTED_35;
        run_test(35, 7);

        test_pixels   = PIXELS_36;
        test_expected = EXPECTED_36;
        run_test(36, 9);

        test_pixels   = PIXELS_37;
        test_expected = EXPECTED_37;
        run_test(37, 7);

        test_pixels   = PIXELS_38;
        test_expected = EXPECTED_38;
        run_test(38, 9);

        test_pixels   = PIXELS_39;
        test_expected = EXPECTED_39;
        run_test(39, 9);

        test_pixels   = PIXELS_40;
        test_expected = EXPECTED_40;
        run_test(40, 8);

        test_pixels   = PIXELS_41;
        test_expected = EXPECTED_41;
        run_test(41, 4);

        test_pixels   = PIXELS_42;
        test_expected = EXPECTED_42;
        run_test(42, 4);

        test_pixels   = PIXELS_43;
        test_expected = EXPECTED_43;
        run_test(43, 2);

        test_pixels   = PIXELS_44;
        test_expected = EXPECTED_44;
        run_test(44, 5);

        test_pixels   = PIXELS_45;
        test_expected = EXPECTED_45;
        run_test(45, 5);

        test_pixels   = PIXELS_46;
        test_expected = EXPECTED_46;
        run_test(46, 4);

        test_pixels   = PIXELS_47;
        test_expected = EXPECTED_47;
        run_test(47, 8);

        test_pixels   = PIXELS_48;
        test_expected = EXPECTED_48;
        run_test(48, 9);

        test_pixels   = PIXELS_49;
        test_expected = EXPECTED_49;
        run_test(49, 6);


        $display("\n====================================================");
        if (errors == 0)
            $display("ALL 50 TESTS PASSED (%0d checks)", total_checks);
        else
            $display("FAILED: %0d errors out of %0d checks", errors, total_checks);
        $display("====================================================\n");
        #50; $finish;
    end

    initial begin #500000000; $display("TIMEOUT"); $finish; end

endmodule
