`timescale 1ns/1ps

module tb_layer_one_digits;

    // ============================================================================
    // Test Parameters - Multiple MNIST-style digits
    // ============================================================================

    // Digit 0
    reg [783:0] TEST_PIXELS_DIGIT_0 = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111110000000000000011110000000111100000000000011110000000001111000000000011110000000000011110000000001110000000000000111000000001111000000000000011110000000111000000000000000111000000011100000000000000011100000001110000000000000001110000000111000000000000000111000000011100000000000000011100000001111000000000000011110000000011100000000000001110000000001111000000000001111000000000011110000000001111000000000000111100000001111000000000000001111111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_OUTPUT_DIGIT_0 = 1568'b11111111111111111111111111111111100001111111100111100111110011111100111100111111101111011111111011110111111110111101111111001111101111110011111001111011111111100001111111111111111111111111111111111111111111111111111111111111111111111111111110110001111111011111101111110111111101111101111111101111011111111011110111111101111101111111011111101111101111111101111111111111111111111111111111111111000000000000000000000000000000000000000000000001111100000010000001100001101000001100010000000010000100000000100001100000001010001100000010100001100000000000001111110000000000000000000000000000000000000000000000000000000000000000011111100000001111111100000111000011100001100000011000111000000110001100000001100011100000011000011100000110000011000011100000111111110000000000010000000000000000001111111111111111111111111111111110000011111110011110011111100111110011111011111110111100111111100111001111111001110011111110111110011111101111110011100011111111111101111111111111111111111111111111000000000000000000000000000000000111111000000011111111000001110000111000011000000110001110000001100011000000011000111000000110000111000001100000110000111000001111111100000000000100000000000000000000000000000000000000000000000000111110000000011000011000001110000111000011000000110000100000000100001000000001000011000000110000111000001100000111001110000000011110000000000000000000000000000000000000000000000000000000000000000001000110000001111111010000111000111010001100000111100111000000110001100000001100011010000011100111110000110000110100011100000111111110000000111110000000000000000000;

    // Digit 1
    reg [783:0] TEST_PIXELS_DIGIT_1 = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111111000000000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_OUTPUT_DIGIT_1 = 1568'b11111111111111111111111111111111000000111111111110011111111111100111111111111001111111111110011111111111100111111111111001111111111110001111111111100111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110111111111111101111111111111011111111111110111111111111101111111111111011111111111110111111111111101111111111111111111111111111111111000000000000000000000000000000001000000000000011110111000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000011000000000000000000000000000000000000000000000000000000000000000000011111110000000111111100000000011100000000000111000000000001110000000000011100000000000111000000000001111000000000011110000000000111000000000000100000000000000000001111111111111111111111111111111110000001111111111001111111111110011111111111100111111111111001111111111110011111111111100111111111111000111111111110001111111111110111111111111111111111111111111111000000000000000000000000000000000111111100000001111111000000000111000000000001110000000000011100000000000111000000000001110000000000011110000000000111100000000001110000000000001000000000000000000000000000000000000000000000000000111111100000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001110000000000011100000000000110000000000000000000000000000000000000000000000000000000000000000000000001000000111111100000000011100000000000111000000000001110000000000011100000000000111000000000001111100000000011110000000000111000000000001100000000000000000000;

    // Digit 2
    reg [783:0] TEST_PIXELS_DIGIT_2 = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000001111111111111111000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111100000000000111100000000001111000000000111100000000000011111000001111100000000000000111111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_OUTPUT_DIGIT_2 = 1568'b11111111111111111111111111111110000000111111111111011111111111101111111111110111111111111011111111111101111111111110111111111111001111111111111001111001111111000000111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111110111111111111011111111111101111111111110111111111111011111111111101111111111111011111111111111011111011111111100011111111111111111111000000000000000000000000000000100000000000001111111011000000000000000000000000000000000000000000000000000000000000000000000001000000000000011000000000000011100010000000011111100000000000000000000000000000000000000000000000001111111110000011111111100000000001110000000000111000000000011100000000001110000000000111000000000011100000010000111100011100000111111110000000111111000000000000000001111111111111111111111111111111000000001111111111100111111111110001111111111000111111111100011111111110001111111111000111111111110011111111111100111100011111100000101111111111111111111111111111111000000000000000000000000000000011111111100000111111111000000000011100000000001110000000000111000000000011100000000001110000000000111000000100001111000111000001111111100000001111110000000000000000000000000000000000000000000000001111111100000000001110000000000011000000000001100000000000110000000000011000000000001100000000000110000000000000110000110000001111111100000000000000000000000000000000000000000000000000000000000000000000001000011111111100000000001110000000000111000000000011100000000001110000000000111000000000011100000001000110110011100001110001110000001111111000000000000000000;

    // Digit 5
    reg [783:0] TEST_PIXELS_DIGIT_5 = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111110000000000000001111100001111110000000000001111000000001111100000000001111000000000011110000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000000000000000000000011110000000000000000000000000111110000000000000000000000000111111111111100000000000000000111111111110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_OUTPUT_DIGIT_5 = 1568'b11111111111111111111111111111111100001111111110011100111111011111100111100111111111111101111111111111001111111111111110000011111111111100111111111111001111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111011001111111101111100111110111111111111101111111111111101111111111111100111111111111111110111111111111101111111111111011111111000000111111111111111111000000000000000000000000000000000000000000000000111100000000010001111000100000000000001100000000000001100000000000001111110000000000000100000000000001000000010000000000000111111111000000000000000000000000000000000000000000000000011111100000001111111110000011100011100001110000001000011100000000000111100001000000111111110000000000001100000000000011000000111111110000001111111100000000000000001111111111111111111111111111111110000011111111001110001111100111111111111001111111111110011111111111110011111111111111111001111111111111011111111111110111111100000001111111111111111111111111111111000000000000000000000000000000000111111000000011111111100000111000111000011100000010000111000000000001111000010000001111111100000000000011000000000000110000001111111100000011111111000000000000000000000000000000000000000000000000011110000000001110111000000110000111000011000000000000111000000000000111000000000000001111100000000000011000000000000110000000111111100000000000000000000000000000000000000000000000000000000000000001000110000000111111011000011100111100001110000111000011110000000000111010000100000111111110000000011111100000000000011000000000001110000001111111100000000000000000;

    // Digit 7
    reg [783:0] TEST_PIXELS_DIGIT_7 = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111111111111111111000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    reg [1567:0] EXPECTED_OUTPUT_DIGIT_7 = 1568'b11111111111111111111111111111111111001111111111110011111111111001111111111110011111111111001111111111110011111111111001111111111110011111111111001111111111100010000011111111111111111111111111111111111111111111111111111111111111111101111111111111011111111111101111111111111011111111111101111111111111011111111111101111111111111011111111111101111111111110011111111111100000000011111111111111111000000000000000000000000000000000001010000000000110100000000001010000000000110100000000001010000000000110100000000001010000000000110100000000001010000000000100000000000001111111111000000000000000000000000000000000000000100000000000011000000000000110000000000011100000000000110000000000011100000000000110000000000011100000000000110000000000011100000000001111111110000011111111100000000000000001111111111111111111111111111111111110111111111111101111111111110111111111111101111111111110111111111111101111111111110111111111111101111111111110111111111111000000001111111111111111111111111111111000000000000000000000001000000000000110000000000001100000000000111000000000001100000000000111000000000001100000000000111000000000001100000000000111000000000011111111100000111111111000000000000000000000000000000000000000000000000000110000000000001100000000000110000000000001100000000000110000000000001100000000000110000000000001100000000000110000000000011111111100000000000000000000000000000000000000000000000000000010000000000011100000000000110000000000011100000000000110000000000011100000000000110000000000011100000000000110000000000011100000000001110000001000011111111100000000000000000;

    // Common weights for all digit tests
    reg [71:0] TEST_WEIGHTS_DIGITS = 72'b111101100000000110101011011111000001011100111111110101110100001000100010;

    // Testbench signals
    reg clk;
    reg rst_n;
    reg [2:0] state;
    reg [783:0] pixels;
    reg [71:0] weights;
    wire [1567:0] layer_one_out;
    wire done;

    // Error tracking
    integer errors = 0;
    integer total_checks = 0;

    // Instantiate DUT
    layer_one dut (
        .clk(clk),
        .rst_n(rst_n),
        .state(state),
        .pixels(pixels),
        .weights(weights),
        .layer_one_out(layer_one_out),
        .done(done)
    );

    // State definitions
    localparam [2:0] s_IDLE    = 3'b000;
    localparam [2:0] s_LOAD    = 3'b001;
    localparam [2:0] s_LAYER_1 = 3'b010;
    localparam [2:0] s_LAYER_2 = 3'b011;
    localparam [2:0] s_LAYER_3 = 3'b100;

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Helper function to get output index
    function integer out_idx;
        input integer w, r, c;
        begin
            out_idx = w*196 + r*14 + c;
        end
    endfunction

    // Verification task
    task verify_output;
        input [1567:0] expected;
        input [7*8:1] digit_name;
        integer w, r, c, idx, mismatches, test_errors;
        begin
            mismatches = 0;
            test_errors = 0;
            $display("\n========================================");
            $display("Verifying Digit %0s Output", digit_name);
            $display("========================================");

            for (w = 0; w < 8; w = w + 1) begin
                for (r = 0; r < 14; r = r + 1) begin
                    for (c = 0; c < 14; c = c + 1) begin
                        idx = out_idx(w, r, c);
                        total_checks = total_checks + 1;

                        if (layer_one_out[idx] !== expected[idx]) begin
                            if (mismatches < 5) begin // Limit error messages
                                $display("ERROR: Mismatch at weight=%0d, row=%0d, col=%0d (idx=%0d)", w, r, c, idx);
                                $display("  Expected: %b, Got: %b",
                                    expected[idx], layer_one_out[idx]);
                            end
                            mismatches = mismatches + 1;
                            test_errors = test_errors + 1;
                        end
                    end
                end
            end

            $display("========================================");
            if (test_errors == 0) begin
                $display("*** DIGIT %0s PASSED ***", digit_name);
                $display("All 1568 outputs match expected values");
            end else begin
                $display("*** DIGIT %0s FAILED ***", digit_name);
                $display("Total errors: %0d / 1568", test_errors);
            end
            $display("========================================\n");

            errors = errors + test_errors;
        end
    endtask

    // Test stimulus
    initial begin
        // Setup VCD dump
        $dumpfile("layer_one.vcd");
        $dumpvars(0, tb_layer_one_digits);

        $display("\n========================================");
        $display("Layer One Testbench - Multiple Digits");
        $display("========================================");
        $display("Testing MNIST-style digits: 0, 1, 2, 5, 7");
        $display("========================================\n");

        errors = 0;
        total_checks = 0;

        // ============================
        // TEST 1: Digit 0
        // ============================
        $display("\n****************************************");
        $display("TEST 1: Digit 0");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_DIGIT_0;
        weights = TEST_WEIGHTS_DIGITS;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_DIGIT_0, "0");

        // ============================
        // TEST 2: Digit 1
        // ============================
        $display("\n****************************************");
        $display("TEST 2: Digit 1");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_DIGIT_1;
        weights = TEST_WEIGHTS_DIGITS;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_DIGIT_1, "1");

        // ============================
        // TEST 3: Digit 2
        // ============================
        $display("\n****************************************");
        $display("TEST 3: Digit 2");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_DIGIT_2;
        weights = TEST_WEIGHTS_DIGITS;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_DIGIT_2, "2");

        // ============================
        // TEST 4: Digit 5
        // ============================
        $display("\n****************************************");
        $display("TEST 4: Digit 5");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_DIGIT_5;
        weights = TEST_WEIGHTS_DIGITS;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_DIGIT_5, "5");

        // ============================
        // TEST 5: Digit 7
        // ============================
        $display("\n****************************************");
        $display("TEST 5: Digit 7");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_DIGIT_7;
        weights = TEST_WEIGHTS_DIGITS;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_DIGIT_7, "7");

        // ============================
        // Final Summary
        // ============================
        $display("\n========================================");
        $display("FINAL TEST SUMMARY");
        $display("========================================");
        if (errors == 0) begin
            $display("*** ALL DIGIT TESTS PASSED ***");
            $display("Tested digits: 0, 1, 2, 5, 7");
            $display("Total checks: %0d", total_checks);
        end else begin
            $display("*** SOME TESTS FAILED ***");
            $display("Total errors: %0d / %0d checks", errors, total_checks);
        end
        $display("========================================\n");

        // End simulation
        #50;
        $finish;
    end

    // Timeout watchdog
    initial begin
        #100000000; // 100ms timeout
        $display("\nERROR: Simulation timeout!");
        $finish;
    end

endmodule
