`timescale 1ns/1ps

module tb_layer_one_simple;

    // ============================================================================
    // Test Parameters - Multiple Test Patterns
    // ============================================================================

    // All Zeros Test
    reg [783:0] TEST_PIXELS_ZEROS = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // All Ones Test
    reg [783:0] TEST_PIXELS_ONES = 784'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

    // MNIST digit '3' - 28x28 flattened to 784 bits
    reg [783:0] TEST_PIXELS_MNIST = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111111110000000000000000111100011111000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000000110000000000000000000000000001100000000000000000000000000111000000000000000000000000000111111000000000000000000000111111100000000000000000000111111110000000000000000001100000000000000000000000000111100000000000000000000011000000000000000000000000011000000000000000000000000001110000000000000000000000000011111111111100000000000000000111111111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Simple weights for all tests - 3x3x8 flattened to 72 bits
    reg [71:0] TEST_WEIGHTS_SIMPLE = 72'b100001111110101010011011001001101111001110000110001111001000000000100000;

    // Weights from Python model (for MNIST test)
    reg [71:0] TEST_WEIGHTS_MNIST = 72'b011000001110000011000000011000011011000111110001000111110001111001010111;

    // Expected outputs
    reg [1567:0] EXPECTED_OUTPUT_ZEROS = 1568'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

    reg [1567:0] EXPECTED_OUTPUT_ONES = 1568'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000111111111111111111111111111110000000000000100000000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000111111111111110000000000000100000000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000010000000000000100000000000001000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111;

    reg [1567:0] EXPECTED_OUTPUT_MNIST = 1568'b00000000000000000000000000000000000110000000001111111000000001100000000000011000000000000010000000000000111100000000011011000000010110000000000110000000000001111111000000000111000000000000000000000000000000000000000000000000000010111110000000111111110000000110000000000001100000000000001100000000000001111000000001111110000001011100000000011000000000000011111110000000001100000000000000000000000000000000000000000000000000000011101000000001101111000000001000000000000010000000000000110000000000000111100000000111001000000000010000000000100000000000001111111000000000010000000000000000000000000000000000000001111110000000111111110000000010000000000001100000000000001110000000000001111000000001111100000001111000000000011000000000000111111110000000001100000000000000000000000000000000001111111111111111111111111111111111100011111111100110011111111101111111111111011111111111111011111111111110001111111111011111111111111111111111110111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111110011001111111111111111111111101111111111111111111111111111100111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111001000111111111011111111111110111111111111100111111111111110001111111111011111111111111111111111011111111111111000000111111111111111111111111111111110000000000000000000111111000000011111111000000010100000000000111000000000000011000000000000111100000000111111000000101110000000001100000000000011111111000000001111000000000000000000000000000000000;
    
    // Testbench signals
    reg clk;
    reg rst_n;
    reg [2:0] state;
    reg [783:0] pixels;
    reg [71:0] weights;
    wire [1567:0] layer_one_out;
    wire done;

    // Error tracking
    integer errors = 0;
    integer total_checks = 0;

    // Instantiate DUT
    layer_one dut (
        .clk(clk),
        .rst_n(rst_n),
        .state(state),
        .pixels(pixels),
        .weights(weights),
        .layer_one_out(layer_one_out),
        .done(done)
    );

    // State definitions
    localparam [2:0] s_IDLE    = 3'b000;
    localparam [2:0] s_LOAD    = 3'b001;
    localparam [2:0] s_LAYER_1 = 3'b010;
    localparam [2:0] s_LAYER_2 = 3'b011;
    localparam [2:0] s_LAYER_3 = 3'b100;

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Helper function to get output index
    function integer out_idx;
        input integer w, r, c;
        begin
            out_idx = w*196 + r*14 + c;
        end
    endfunction

    // Verification task
    task verify_output;
        input [1567:0] expected;
        integer w, r, c, idx, mismatches, test_errors;
        begin
            mismatches = 0;
            test_errors = 0;
            $display("\n========================================");
            $display("Verifying Output Against Python Model");
            $display("========================================");

            for (w = 0; w < 8; w = w + 1) begin
                for (r = 0; r < 14; r = r + 1) begin
                    for (c = 0; c < 14; c = c + 1) begin
                        idx = out_idx(w, r, c);
                        total_checks = total_checks + 1;

                        if (layer_one_out[idx] !== expected[idx]) begin
                            if (mismatches < 10) begin // Limit error messages
                                $display("ERROR: Mismatch at weight=%0d, row=%0d, col=%0d (idx=%0d)", w, r, c, idx);
                                $display("  Expected: %b, Got: %b",
                                    expected[idx], layer_one_out[idx]);
                            end
                            mismatches = mismatches + 1;
                            test_errors = test_errors + 1;
                        end
                    end
                end
                if (mismatches == 0) begin
                    $display("Weight %0d: PASS (all 196 outputs correct)", w);
                end else begin
                    $display("Weight %0d: %0d mismatches", w, mismatches);
                end
            end

            $display("========================================");
            if (test_errors == 0) begin
                $display("*** TEST PASSED ***");
                $display("All 1568 outputs match expected values");
            end else begin
                $display("*** TEST FAILED ***");
                $display("Total errors in this test: %0d / 1568", test_errors);
            end
            $display("========================================\n");

            errors = errors + test_errors;
        end
    endtask

    // Test stimulus
    initial begin
        $display("\n========================================");
        $display("Layer One Testbench - Multiple Tests");
        $display("========================================");
        $display("Running 3 test cases:");
        $display("  1. All zeros");
        $display("  2. All ones");
        $display("  3. MNIST digit '3'");
        $display("========================================\n");

        errors = 0;
        total_checks = 0;

        // ============================
        // TEST 1: All Zeros
        // ============================
        $display("\n****************************************");
        $display("TEST 1: All Zeros Pattern");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_ZEROS;
        weights = TEST_WEIGHTS_SIMPLE;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete (done asserted)", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_ZEROS);

        // ============================
        // TEST 2: All Ones
        // ============================
        $display("\n****************************************");
        $display("TEST 2: All Ones Pattern");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_ONES;
        weights = TEST_WEIGHTS_SIMPLE;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete (done asserted)", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_ONES);

        // ============================
        // TEST 3: MNIST Digit '3'
        // ============================
        $display("\n****************************************");
        $display("TEST 3: MNIST Digit '3'");
        $display("****************************************");

        rst_n = 0;
        state = s_IDLE;
        pixels = TEST_PIXELS_MNIST;
        weights = TEST_WEIGHTS_MNIST;

        #20;
        rst_n = 1;
        $display("[%0t] Reset released", $time);

        #20;
        state = s_LAYER_1;
        $display("[%0t] Starting LAYER_1 processing", $time);

        wait(done == 1);
        $display("[%0t] Processing complete (done asserted)", $time);
        #100;

        verify_output(EXPECTED_OUTPUT_MNIST);

        // ============================
        // Final Summary
        // ============================
        $display("\n========================================");
        $display("FINAL TEST SUMMARY");
        $display("========================================");
        if (errors == 0) begin
            $display("*** ALL TESTS PASSED ***");
            $display("Total checks: %0d", total_checks);
        end else begin
            $display("*** SOME TESTS FAILED ***");
            $display("Total errors: %0d / %0d checks", errors, total_checks);
        end
        $display("========================================\n");

        // End simulation
        #50;
        $finish;
    end

    // Waveform dumping
    initial begin
        $dumpfile("layer_one.vcd");
        $dumpvars(0, tb_layer_one_simple);
    end

    // Timeout watchdog
    initial begin
        #500000;
        $display("\n========================================");
        $display("ERROR: Simulation timeout!");
        $display("========================================");
        $finish;
    end

endmodule
